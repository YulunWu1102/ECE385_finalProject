module rtank_rom ( input [15:0]	addr,
						 input [1:0] tankSelection,
						output [3:0]	data
					 );

	parameter ADDR_WIDTH = 16;
   parameter DATA_WIDTH =  4;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:3499][3:0] R_ROM = {


4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0
// above are rtank



        };
		  
		  
		  
parameter [0:3499][3:0] G_ROM = {


4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h4,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h5,
4'h4,
4'h4,
4'h4,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h5,
4'h4,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h5,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h5,
4'h4,
4'h4,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h4,
4'h4,
4'h4,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,

// above are gtank



        };
		  
		  
parameter [0:3499][DATA_WIDTH-1:0] B_ROM = {

4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h9,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h9,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h9,
4'h9,
4'h7,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h8,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h7,
4'h7,
4'h7,
4'h8,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h9,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h8,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h8,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h8,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h8,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h8,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h8,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h8,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h8,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h8,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h8,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h9,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h8,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h7,
4'h7,
4'h7,
4'h7,
4'h7,
4'h8,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h9,
4'h9,
4'h7,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h8,
4'h7,
4'h7,
4'h7,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h7,
4'h7,
4'h7,
4'h8,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,

// above are btank



        };

		  
		  
	always_comb begin:tank_select
	
	case(tankSelection)
	
	2'b00: begin
		data = R_ROM[addr];
	
	end
	
	2'b01: begin
		data = G_ROM[addr];	
	end
	
	2'b10: begin
		data = B_ROM[addr];
	end
	
	2'b11: begin
		data = B_ROM[addr];
	end
	
	default:;
	
	endcase
	
	end



endmodule  