module num_rom ( input [12:0]	addr,
						 input [3:0] currNum,
						output [3:0]	data
					 );

	// ROM definition
	// numx: x from 0 to 9
	// each number is 20 x 30 (width x height)
	// selection logic missing

		
	parameter [0:599][3:0] num0 = {
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hc,
4'h3,
4'hd,
4'h3,
4'h3,
4'hc,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h3,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h3,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'h3,
4'h6,
4'h6,
4'h6,
4'h6,
4'h3,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hc,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'h2,
4'h2,
4'h2,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1
	};

	parameter [0:599][3:0] num1 = {
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'hf,
4'h6,
4'h6,
4'hf,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1
	};

	parameter [0:599][3:0] num2 = {
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'hc,
4'h3,
4'h2,
4'h2,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'h3,
4'h3,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h6,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h6,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h3,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'hc,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'hd,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'h4,
4'h6,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'h3,
4'hc,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'hc,
4'h3,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1
	};

	parameter [0:599][3:0] num3 = {
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'hc,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'h3,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'hd,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'h2,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'hd,
4'hc,
4'h3,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h3,
4'h4,
4'h6,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'h3,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'h3,
4'hf,
4'hf,
4'hf,
4'hf,
4'h3,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hc,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1
	};

	parameter [0:599][3:0] num4 = {
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h3,
4'h4,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h4,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'h2,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h6,
4'h3,
4'h3,
4'h6,
4'h3,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hc,
4'hc,
4'hc,
4'hc,
4'hc,
4'hc,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1
	};

	parameter [0:599][3:0] num5 = {
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h3,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'h6,
4'hf,
4'hf,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hc,
4'h2,
4'h2,
4'h2,
4'hc,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'hc,
4'h2,
4'h2,
4'he,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'h3,
4'h6,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h3,
4'hd,
4'hd,
4'h3,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1
	};

	parameter [0:599][3:0] num6 = {
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hc,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h3,
4'hd,
4'hd,
4'h3,
4'h2,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h3,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'h3,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'hf,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h6,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h2,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'hc,
4'h1,
4'h1,
4'h2,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'he,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'hc,
4'h1,
4'h1,
4'h2,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'hc,
4'h1,
4'h1,
4'h2,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h3,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hc,
4'hd,
4'hd,
4'h3,
4'h3,
4'h3,
4'h3,
4'hd,
4'hd,
4'h3,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'he,
4'he,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1
	};

	parameter [0:599][3:0] num7 = {
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'he,
4'he,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1
	};

	parameter [0:599][3:0] num8 = {
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'hf,
4'h3,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hf,
4'h4,
4'h4,
4'hf,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'h6,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h3,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'h2,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h2,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'he,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h2,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'hc,
4'he,
4'hc,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'h3,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h3,
4'hd,
4'h3,
4'h6,
4'h4,
4'h4,
4'h4,
4'hf,
4'h3,
4'hd,
4'h3,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'hd,
4'hd,
4'hd,
4'h3,
4'h3,
4'hd,
4'hd,
4'h2,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1
	};

	parameter [0:599][3:0] num9 = {
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'h3,
4'h6,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'h1,
4'h1,
4'h2,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h3,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h3,
4'h4,
4'h6,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h3,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h6,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h3,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h3,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'h6,
4'h4,
4'h4,
4'h4,
4'hf,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'h3,
4'hd,
4'hd,
4'h3,
4'h6,
4'h3,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hc,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'hc,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1
	};

		    
 always_comb begin:num_select
 
 case(currNum)
 
 0: begin
  data = num9[addr];
  end
 
 1: begin
  data = num8[addr];
  end
  
  2: begin
  data = num7[addr];
  end
 3: begin
  data = num6[addr];
  end
  
  4: begin
  data = num5[addr];
  end
  
  5: begin
  data = num4[addr];
  end
  
  6: begin
  data = num3[addr];
  end
  
  7: begin
  data = num2[addr];
  end
  
   8: begin
  data = num1[addr];
  end
 
   9: begin
  data = num0[addr];
  end
  
  9: begin
  data = num0[addr];
  end
  
  10: begin
  data = num0[addr];
  end
  
  11: begin
  data = num0[addr];
  end
  
  12: begin
  data = num0[addr];
  end
  
  13: begin
  data = num0[addr];
  end
  
  14: begin
  data = num0[addr];
  end
  
  15: begin
  data = num0[addr];
  end
  

 default:;
 
 endcase
 
 end

 endmodule

