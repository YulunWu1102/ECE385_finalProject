module font_rom ( input [15:0]	addr,
						output [7:0]	data
					 );

	parameter ADDR_WIDTH = 11;
   parameter DATA_WIDTH =  8;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:3499][DATA_WIDTH-1:0] ROM = {
       8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000010,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000001,
8'b00000001,
8'b00000001,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000
// above are rtank

        };

	assign data = ROM[addr];

endmodule  