module bullet_rom ( input [13:0]	addr,
						 input [1:0] tankSelection,					 
						 output [3:0]	data
					 );


				
	// ROM definition
	// BU1, BU2, BU3	
	// missing selection logic in the end

		

	parameter [0:399][3:0] BU0 = {
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h4,
4'h7,
4'h7,
4'hb,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h7,
4'h1,
4'h7,
4'h2,
4'h0,
4'h0,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'hb,
4'hb,
4'hc,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h8,
4'ha,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h8,
4'h8,
4'h8,
4'h9,
4'h9,
4'hd,
4'h9,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h8,
4'h8,
4'he,
4'h8,
4'h8,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h8,
4'he,
4'he,
4'he,
4'h8,
4'h8,
4'h9,
4'h9,
4'ha,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h8,
4'he,
4'he,
4'he,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h9,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h9,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h9,
4'h9,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h9,
4'h8,
4'h8,
4'h8,
4'h8,
4'h8,
4'h9,
4'h9,
4'h8,
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'h9,
4'h8,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h9,
4'h9,
4'h9,
4'h9,
4'h9,
4'ha,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0

	};

	parameter [0:399][3:0] BU1 = {
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'h0,
4'h2,
4'h2,
4'h7,
4'h7,
4'h4,
4'h7,
4'h7,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h4,
4'h7,
4'h7,
4'h7,
4'he,
4'h7,
4'h4,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h0,
4'h0,
4'h2,
4'h6,
4'hf,
4'hf,
4'hf,
4'h4,
4'h7,
4'h7,
4'he,
4'he,
4'h1,
4'hb,
4'hf,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'hf,
4'hf,
4'hf,
4'hb,
4'h7,
4'h1,
4'he,
4'he,
4'h1,
4'h4,
4'hf,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h4,
4'h2,
4'hf,
4'h4,
4'hf,
4'hf,
4'hf,
4'h4,
4'h7,
4'he,
4'h1,
4'h1,
4'h1,
4'h4,
4'hf,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h4,
4'h4,
4'hf,
4'hf,
4'h4,
4'h7,
4'h7,
4'he,
4'h1,
4'he,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'hf,
4'h2,
4'h2,
4'h2,
4'hf,
4'hf,
4'hf,
4'hb,
4'h7,
4'h7,
4'h7,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'hf,
4'h4,
4'h4,
4'hf,
4'hf,
4'hf,
4'hf,
4'h4,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'hf,
4'hf,
4'hf,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h4,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0

	};

	parameter [0:399][3:0] BU2 = {
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'hc,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'hc,
4'h2,
4'h2,
4'h2,
4'h2,
4'hc,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'hc,
4'hc,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'hc,
4'hc,
4'h2,
4'hc,
4'hc,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'hc,
4'hc,
4'hc,
4'hc,
4'hc,
4'hc,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'hc,
4'hc,
4'hc,
4'h3,
4'hc,
4'h2,
4'hc,
4'hc,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'hc,
4'hc,
4'hc,
4'h3,
4'hc,
4'h2,
4'hc,
4'hc,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'hc,
4'hc,
4'hc,
4'hc,
4'h3,
4'h3,
4'h3,
4'hc,
4'hc,
4'hc,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'hc,
4'hc,
4'hc,
4'hc,
4'hc,
4'hc,
4'h3,
4'h3,
4'h3,
4'h3,
4'hc,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'hc,
4'hc,
4'hc,
4'h2,
4'h2,
4'hc,
4'hc,
4'hc,
4'hc,
4'h3,
4'h3,
4'h3,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'hc,
4'hb,
4'h2,
4'h2,
4'he,
4'h2,
4'hc,
4'hc,
4'hc,
4'hc,
4'h3,
4'h3,
4'hc,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'hc,
4'hc,
4'hc,
4'h2,
4'h2,
4'hc,
4'hc,
4'hc,
4'hc,
4'hc,
4'h3,
4'hd,
4'hc,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'hc,
4'hc,
4'hc,
4'h2,
4'h2,
4'hc,
4'hc,
4'hc,
4'h3,
4'h3,
4'hd,
4'h3,
4'hc,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'hc,
4'hc,
4'hc,
4'hc,
4'hc,
4'hc,
4'hc,
4'hc,
4'hc,
4'h3,
4'hd,
4'h3,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'hc,
4'hc,
4'hc,
4'hc,
4'hc,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'hd,
4'h3,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'hc,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'hd,
4'h3,
4'hc,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'hd,
4'hd,
4'h3,
4'h0,
4'h2,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h3,
4'hd,
4'h3,
4'h3,
4'h2,
4'h0,
4'h0,
4'h2,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0

	};
	
	 always_comb begin:bullet_select
	 
		 case(tankSelection)
		 
			 2'b00: begin
				data = BU0[addr];
			 
			 end
			 
			 2'b01: begin
				data = BU1[addr]; 
			 end
			 
			 2'b10: begin
				data = BU2[addr];
			 end
			 
			 2'b11: begin
				data = BU2[addr];
			 end
			 
			 default:;
		 
		 endcase
	 
	 end

 endmodule
 