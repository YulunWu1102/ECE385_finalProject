module hp_rom ( input [13:0]	addr,
					 input [3:0] HPSelection,
					 output [7:0]	data
					 );

	// ROM definition
	// 11 different states of HP
	// HPx, x goes from 10 to 0 
	// HPSelection logic not implemented

		
	parameter [0:1399][7:0] HP10 = {
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h21,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h61,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01


	};


	parameter [0:1399][7:0] HP9 = {
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h21,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h61,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01


	};

	parameter [0:1399][7:0] HP8 = {
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h21,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h61,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01


	};


	parameter [0:1399][7:0] HP7 = {
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h21,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h61,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01


	};

	parameter [0:1399][7:0] HP6 = {
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h21,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h61,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01


	};

	parameter [0:1399][7:0] HP5 = {
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h21,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h61,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01


	};

	parameter [0:1399][7:0] HP4 = {
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h21,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h61,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01


	};

	parameter [0:1399][7:0] HP3 = {
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h21,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h61,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01


	};

	parameter [0:1399][7:0] HP2 = {
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h41,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h21,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h61,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01


	};

	parameter [0:1399][7:0] HP1 = {
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'hf1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h21,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h61,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01


	};

	parameter [0:1399][7:0] HP0 = {
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h21,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h61,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h61,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'hd1,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01,
8'h01

	};
	
always_comb begin:hp_func
	 
		 case(HPSelection)
		 
			 0: data = HP0[addr];
			 1: data = HP1[addr];
			 2: data = HP2[addr];
			 3: data = HP3[addr];
			 4: data = HP4[addr];
			 5: data = HP5[addr];
			 6: data = HP6[addr];
			 7: data = HP7[addr];
			 8: data = HP8[addr];
			 9: data = HP9[addr];
			 10: data = HP10[addr];
			 
			 default: data = HP10[addr];
		 
		 endcase
	 
	 end

 endmodule
 
