module background_rom ( input [18:0]	addr,
						output [3:0]	data
					 );

	//parameter ADDR_WIDTH = 19;
   //parameter DATA_WIDTH =  4;
	//logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:38399][4:0] ROM = {

4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'hb,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'h5,
4'hb,
4'h5,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h0,
4'ha,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'h5,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'hb,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'h0,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'hb,
4'h6,
4'h6,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h0,
4'h0,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h0,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h5,
4'h5,
4'h5,
4'h5,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h0,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h0,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h0,
4'h0,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h0,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h0,
4'h0,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'ha,
4'ha,
4'ha,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'hb,
4'hb,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'h6,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h0,
4'h0,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h0,
4'h6,
4'h6,
4'h6,
4'h6,
4'hb,
4'hb,
4'h4,
4'h4,
4'hb,
4'h6,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'ha,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h6,
4'h6,
4'hb,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h5,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h5,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'hb,
4'hb,
4'hb,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'hb,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h0,
4'h0,
4'h6,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'hb,
4'hb,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'hb,
4'h4,
4'h4,
4'h4,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'hb,
4'hb,
4'hb,
4'h4,
4'h0,
4'h0,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h0,
4'h6,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h6,
4'h6,
4'h0,
4'h0,
4'h0,
4'h0,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hd,
4'hd,
4'h4,
4'h4,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'hb,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'hb,
4'hb,
4'hb,
4'hb,
4'h0,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h0,
4'h0,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'h0,
4'h0,
4'h0,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'h0,
4'h0,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'hb,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'h0,
4'h0,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h0,
4'h0,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'hb,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'h1,
4'h1,
4'h1,
4'hf,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'h1,
4'h1,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'h1,
4'h1,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'h1,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'hd,
4'hd,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'hf,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'hf,
4'hf,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'hf,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hf,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hf,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hf,
4'hf,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hf,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'he,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1



        };

	assign data = ROM[addr];

endmodule  