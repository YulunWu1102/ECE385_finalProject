module rtank_rom ( input [15:0]	addr,
						 input [1:0] tankSelection, Direction,						 
						 output [7:0]	data
					 );

	parameter ADDR_WIDTH = 16;
   parameter DATA_WIDTH =  4;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition
	// 三个坦克是 R， Y(之前是G)， B . R_ROM_X: X = left or right	 (X is L or R)	
	// 4/26 add four explosion 50x50 each. Name: EXP1, EXP2, EXP3, EXP4
	// added 8'hAB, A is the color pallette number, B is the priority number (6 is highest, 0 is lowest)
	// Priority: 6: explosion; 5: tank2; 4: tank1; 3: bullet; 2: 血条2; 1: 血条1; 0: Background 
	// deleted selection at the end

		

	parameter [0:6999][7:0] R_ROM = {
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h25,
8'h65,
8'h65,
8'hf5,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h65,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h65,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'h65,
8'hf5,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h35,
8'h35,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h35,
8'h25,
8'h25,
8'hc5,
8'hc5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h25,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hc5,
8'h25,
8'h35,
8'hf5,
8'h35,
8'hd5,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h65,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h65,
8'h35,
8'hc5,
8'hc5,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'hc5,
8'h25,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'hf5,
8'h45,
8'hf5,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'hf5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'hc5,
8'hd5,
8'h65,
8'h45,
8'hf5,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h65,
8'h65,
8'hf5,
8'hf5,
8'h65,
8'h65,
8'h65,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h65,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hc5,
8'hc5,
8'h35,
8'h65,
8'h45,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h65,
8'h65,
8'h35,
8'h65,
8'h65,
8'hf5,
8'hf5,
8'h65,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'hd5,
8'h45,
8'h45,
8'hf5,
8'hf5,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h35,
8'h65,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'h35,
8'h35,
8'h65,
8'h65,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h45,
8'h45,
8'hf5,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'hf5,
8'h65,
8'h65,
8'h65,
8'h65,
8'h35,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hc5,
8'h45,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h65,
8'hf5,
8'h65,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h65,
8'h45,
8'hf5,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h65,
8'hf5,
8'hf5,
8'h65,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'hf5,
8'h65,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'hf5,
8'h65,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h35,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'hf5,
8'h65,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h35,
8'h65,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h65,
8'h65,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h25,
8'h25,
8'h45,
8'h25,
8'h25,
8'h65,
8'h65,
8'h65,
8'h65,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h65,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h25,
8'h45,
8'hf5,
8'hf5,
8'h45,
8'hf5,
8'h65,
8'hf5,
8'hf5,
8'h65,
8'h65,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h65,
8'h45,
8'h45,
8'hf5,
8'h65,
8'h65,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h65,
8'h65,
8'hf5,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h65,
8'h45,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h45,
8'h45,
8'hf5,
8'h35,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h65,
8'h25,
8'h25,
8'h45,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h45,
8'hf5,
8'hf5,
8'hf5,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h45,
8'h45,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h45,
8'h65,
8'h35,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h25,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h45,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h45,
8'hf5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'hf5,
8'h65,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h35,
8'h65,
8'h65,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h65,
8'hf5,
8'hf5,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h45,
8'h35,
8'hd5,
8'h35,
8'hd5,
8'h35,
8'hf5,
8'h65,
8'hf5,
8'hf5,
8'hf5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hf5,
8'hf5,
8'h65,
8'h65,
8'h35,
8'hd5,
8'h65,
8'h65,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h65,
8'h45,
8'hf5,
8'hf5,
8'hd5,
8'hd5,
8'h35,
8'hd5,
8'h35,
8'hf5,
8'h35,
8'hd5,
8'h35,
8'hd5,
8'h35,
8'hf5,
8'h65,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h65,
8'hf5,
8'hf5,
8'h65,
8'h65,
8'hd5,
8'hd5,
8'h65,
8'h65,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h35,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h35,
8'hf5,
8'h45,
8'hf5,
8'hf5,
8'hf5,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h65,
8'hf5,
8'hd5,
8'hd5,
8'hd5,
8'h65,
8'h65,
8'h65,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h35,
8'h35,
8'hd5,
8'h65,
8'h35,
8'hd5,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'h65,
8'h65,
8'h65,
8'h65,
8'hf5,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h65,
8'h65,
8'h45,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hf5,
8'h65,
8'h65,
8'hf5,
8'hf5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'hf5,
8'h65,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h65,
8'h45,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'h65,
8'h65,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h35,
8'h45,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h35,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h25,
8'h45,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'h35,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h35,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h45,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'hf5,
8'hf5,
8'h65,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h65,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'h25,
8'h65,
8'h65,
8'hf5,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h35,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h65,
8'h65,
8'h65,
8'h25,
8'h05,
8'h05,
8'hd5,
8'h65,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h35,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h65,
8'h65,
8'h65,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'hf5,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'hf5,
8'hf5,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h35,
8'h65,
8'h05,
8'h05,
8'h05,
8'h35,
8'h65,
8'h35,
8'hd5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'hf5,
8'h65,
8'h05,
8'h05,
8'h05,
8'h25,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h65,
8'h35,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h65,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h65,
8'h65,
8'h65,
8'hd5,
8'h65,
8'h65,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'hf4,
8'h64,
8'h64,
8'h24,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'hf4,
8'h64,
8'h64,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'h34,
8'h34,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hc4,
8'hc4,
8'h64,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'hd4,
8'h34,
8'hf4,
8'h34,
8'h24,
8'hc4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'hf4,
8'hf4,
8'h44,
8'hf4,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'h24,
8'hc4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'hc4,
8'hc4,
8'h34,
8'h64,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h64,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'hf4,
8'hf4,
8'h44,
8'h64,
8'hd4,
8'hc4,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hf4,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'h64,
8'hf4,
8'hf4,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'hf4,
8'hf4,
8'hf4,
8'h44,
8'h64,
8'h64,
8'hc4,
8'hc4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h64,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'hf4,
8'h44,
8'h44,
8'hd4,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h24,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h34,
8'h64,
8'h64,
8'h64,
8'h64,
8'hf4,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'hf4,
8'hf4,
8'h44,
8'h44,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h64,
8'h64,
8'h34,
8'h34,
8'hd4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'h64,
8'hf4,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'hf4,
8'hf4,
8'h44,
8'hc4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'h64,
8'hf4,
8'hf4,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'hf4,
8'h44,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h64,
8'hf4,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h34,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'hf4,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h64,
8'h64,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'h34,
8'hd4,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'h04,
8'h04,
8'h64,
8'hc4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'h64,
8'h64,
8'h24,
8'h24,
8'h44,
8'h24,
8'h24,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h64,
8'h64,
8'hf4,
8'h64,
8'hf4,
8'h44,
8'hf4,
8'hf4,
8'h44,
8'h24,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'hd4,
8'hd4,
8'h64,
8'hf4,
8'hf4,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h64,
8'h64,
8'h44,
8'h44,
8'h64,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'hf4,
8'h44,
8'h44,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'h44,
8'h44,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'hf4,
8'hf4,
8'hf4,
8'h44,
8'hc4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'h44,
8'h44,
8'h24,
8'h64,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h64,
8'h64,
8'h64,
8'h64,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'h34,
8'h64,
8'h44,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'hf4,
8'h44,
8'h44,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h34,
8'h64,
8'h64,
8'h64,
8'hf4,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'hf4,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hf4,
8'h44,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'hf4,
8'h44,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'h64,
8'h64,
8'hd4,
8'h34,
8'h64,
8'h64,
8'hf4,
8'hf4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'hf4,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h44,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hf4,
8'hf4,
8'h64,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h34,
8'h64,
8'h64,
8'h64,
8'h64,
8'hd4,
8'hd4,
8'h64,
8'h64,
8'hd4,
8'hd4,
8'h64,
8'h64,
8'hf4,
8'hf4,
8'h64,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'hf4,
8'h34,
8'hd4,
8'h34,
8'hd4,
8'h64,
8'hf4,
8'h34,
8'hd4,
8'h34,
8'hd4,
8'hd4,
8'hf4,
8'hf4,
8'h44,
8'h64,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'hf4,
8'h64,
8'h64,
8'h64,
8'h64,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h34,
8'h34,
8'h64,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'h64,
8'hf4,
8'hd4,
8'hd4,
8'hd4,
8'hf4,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'h44,
8'hf4,
8'h34,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'h34,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'hf4,
8'hf4,
8'h64,
8'hf4,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'h44,
8'h64,
8'h64,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h24,
8'h24,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'h64,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'h44,
8'h64,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h34,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'h44,
8'h34,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h34,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'hd4,
8'hd4,
8'h34,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'h44,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h64,
8'hf4,
8'hf4,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'h44,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h34,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'hf4,
8'hf4,
8'h64,
8'h64,
8'h04,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h34,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'h34,
8'h34,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'h24,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'h34,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h34,
8'h34,
8'hd4,
8'h04,
8'h04,
8'h04,
8'h24,
8'h34,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'hf4,
8'h64,
8'h64,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'h34,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h64,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h64,
8'h64,
8'h64,
8'h64,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04

	};


	
	parameter [0:6999][7:0] Y_ROM = {
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h25,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h95,
8'h95,
8'hd5,
8'hd5,
8'hd5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'he5,
8'he5,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h95,
8'h95,
8'h95,
8'h25,
8'hb5,
8'hb5,
8'h25,
8'h25,
8'ha5,
8'h95,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'ha5,
8'h95,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h25,
8'hb5,
8'h75,
8'h75,
8'h75,
8'hb5,
8'h25,
8'h85,
8'h95,
8'h95,
8'h95,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h25,
8'h75,
8'h75,
8'h75,
8'hb5,
8'h25,
8'h85,
8'h85,
8'h85,
8'h85,
8'h95,
8'h95,
8'h95,
8'h95,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h95,
8'h25,
8'h75,
8'h75,
8'hb5,
8'hc5,
8'h25,
8'hb5,
8'hb5,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'h95,
8'he5,
8'h85,
8'h85,
8'h85,
8'h85,
8'h25,
8'hb5,
8'h75,
8'h75,
8'h75,
8'hb5,
8'h25,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h95,
8'h95,
8'h95,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h85,
8'h75,
8'h75,
8'h75,
8'h75,
8'hc5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'h35,
8'h85,
8'he5,
8'h85,
8'h85,
8'h25,
8'hb5,
8'h75,
8'h75,
8'h75,
8'h75,
8'h25,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h95,
8'ha5,
8'h35,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h25,
8'ha5,
8'he5,
8'h85,
8'h95,
8'hb5,
8'h75,
8'h75,
8'h75,
8'h75,
8'h25,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h95,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h25,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h85,
8'h25,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h25,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h95,
8'h85,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'hb5,
8'h75,
8'h75,
8'h75,
8'h75,
8'hb5,
8'h95,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h85,
8'h85,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hc5,
8'h25,
8'hc5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'ha5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'ha5,
8'ha5,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h25,
8'h05,
8'h05,
8'h25,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h25,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h35,
8'ha5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h25,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'h85,
8'h85,
8'h85,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h25,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h85,
8'h85,
8'h85,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'hd5,
8'hd5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'ha5,
8'h95,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h85,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h35,
8'h25,
8'h25,
8'h25,
8'h25,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'h25,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h25,
8'h25,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'h25,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hc5,
8'hd5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h25,
8'hb5,
8'h75,
8'h75,
8'h25,
8'h25,
8'h25,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'hb5,
8'hb5,
8'h25,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h95,
8'h95,
8'h95,
8'ha5,
8'hc5,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'h25,
8'h25,
8'h25,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'ha5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'ha5,
8'h95,
8'ha5,
8'h95,
8'h95,
8'h25,
8'h25,
8'h25,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'ha5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h25,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'h25,
8'hb5,
8'hb5,
8'hc5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hb5,
8'hc5,
8'ha5,
8'ha5,
8'h95,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'h95,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h25,
8'h25,
8'hb5,
8'hb5,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'hb5,
8'hb5,
8'hb5,
8'h25,
8'h25,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'ha5,
8'ha5,
8'ha5,
8'hc5,
8'hc5,
8'hb5,
8'h25,
8'ha5,
8'h95,
8'ha5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'ha5,
8'h95,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h25,
8'h25,
8'h25,
8'hb5,
8'hb5,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'hb5,
8'hb5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'ha5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'h95,
8'h95,
8'h95,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h25,
8'h25,
8'h25,
8'hb5,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'h75,
8'hb5,
8'hb5,
8'h25,
8'h25,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'hb5,
8'h75,
8'h75,
8'h75,
8'h75,
8'hb5,
8'h25,
8'h25,
8'h25,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'hd5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h25,
8'h25,
8'hb5,
8'hb5,
8'h25,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h25,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'hd4,
8'hd4,
8'hd4,
8'h94,
8'h94,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'h94,
8'h94,
8'h24,
8'h24,
8'h24,
8'hb4,
8'h24,
8'h94,
8'h94,
8'h94,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'he4,
8'he4,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h84,
8'h24,
8'hb4,
8'h74,
8'h74,
8'h74,
8'hb4,
8'h24,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h94,
8'h84,
8'h84,
8'h94,
8'ha4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h84,
8'h84,
8'h84,
8'h84,
8'h24,
8'h74,
8'h74,
8'h74,
8'h74,
8'h24,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h94,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h24,
8'hb4,
8'h74,
8'h74,
8'h74,
8'hb4,
8'h24,
8'h84,
8'h84,
8'h84,
8'h84,
8'he4,
8'h94,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'hb4,
8'hb4,
8'h24,
8'h24,
8'h24,
8'hc4,
8'hb4,
8'h74,
8'h74,
8'h24,
8'h94,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h24,
8'h74,
8'h74,
8'h74,
8'h74,
8'hb4,
8'h84,
8'h84,
8'h84,
8'he4,
8'h84,
8'h34,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'h74,
8'hb4,
8'hb4,
8'hc4,
8'h74,
8'h74,
8'h74,
8'hb4,
8'h84,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'ha4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'hb4,
8'h74,
8'h74,
8'h74,
8'h74,
8'h24,
8'h84,
8'h84,
8'h84,
8'hd4,
8'h24,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'hc4,
8'hc4,
8'h94,
8'h94,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h84,
8'h94,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h24,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h24,
8'h84,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h24,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h84,
8'h84,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h94,
8'hb4,
8'h74,
8'h74,
8'h74,
8'h74,
8'hb4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'ha4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'hc4,
8'h24,
8'h24,
8'hc4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'hd4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'h24,
8'h04,
8'h04,
8'h24,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'h04,
8'h04,
8'h24,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'ha4,
8'h34,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'h24,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h84,
8'h84,
8'h84,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h84,
8'h84,
8'h84,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'h94,
8'ha4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h24,
8'h24,
8'h24,
8'h24,
8'h34,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h84,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'h94,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'hd4,
8'h24,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'h24,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h24,
8'h24,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'h24,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'h24,
8'hb4,
8'hb4,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'h24,
8'h24,
8'h24,
8'h74,
8'h74,
8'hb4,
8'h24,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'ha4,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h24,
8'h24,
8'h24,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'ha4,
8'h94,
8'h94,
8'h94,
8'ha4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'ha4,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'h24,
8'h24,
8'h84,
8'h94,
8'h94,
8'ha4,
8'h94,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'h34,
8'hc4,
8'hb4,
8'hb4,
8'h24,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h24,
8'h94,
8'h94,
8'h94,
8'ha4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h94,
8'ha4,
8'ha4,
8'hc4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'hb4,
8'h24,
8'hb4,
8'hb4,
8'h24,
8'h24,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'h94,
8'ha4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'ha4,
8'h94,
8'ha4,
8'h24,
8'hb4,
8'hc4,
8'hc4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'hc4,
8'hc4,
8'hc4,
8'h24,
8'h24,
8'hb4,
8'hb4,
8'hb4,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'hb4,
8'hb4,
8'h24,
8'h24,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'ha4,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h24,
8'h24,
8'h24,
8'h24,
8'hb4,
8'hb4,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'hb4,
8'hb4,
8'hb4,
8'h24,
8'h24,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'h94,
8'ha4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h24,
8'h24,
8'hb4,
8'hb4,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'h74,
8'hb4,
8'h24,
8'h24,
8'h24,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'h94,
8'h94,
8'ha4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h24,
8'h24,
8'h24,
8'hb4,
8'h74,
8'h74,
8'h74,
8'h74,
8'hb4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'h24,
8'hb4,
8'hb4,
8'h24,
8'h24,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'hd4,
8'hd4,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h24,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04


	};





	parameter [0:6999][7:0] B_ROM = {
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'he5,
8'he5,
8'h25,
8'hc5,
8'h25,
8'h25,
8'h35,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'he5,
8'h15,
8'h15,
8'h25,
8'hc5,
8'h25,
8'h25,
8'h25,
8'h35,
8'hc5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'he5,
8'h15,
8'h15,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'he5,
8'h15,
8'h15,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h25,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'he5,
8'h15,
8'h15,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h25,
8'h25,
8'h25,
8'h25,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'he5,
8'he5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'hd5,
8'h35,
8'h65,
8'h65,
8'h65,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'he5,
8'hc5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hc5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'he5,
8'he5,
8'h25,
8'h35,
8'hc5,
8'hc5,
8'h35,
8'h65,
8'h45,
8'hf5,
8'h65,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h25,
8'h05,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hd5,
8'h35,
8'h35,
8'hc5,
8'h35,
8'h35,
8'h65,
8'h45,
8'h45,
8'h65,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h35,
8'hd5,
8'h35,
8'h35,
8'h35,
8'hc5,
8'hc5,
8'h35,
8'h35,
8'h65,
8'h45,
8'h45,
8'h35,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h05,
8'h05,
8'h25,
8'hd5,
8'ha5,
8'ha5,
8'ha5,
8'hd5,
8'hd5,
8'hc5,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'h35,
8'h35,
8'hd5,
8'h35,
8'h35,
8'h35,
8'hc5,
8'hc5,
8'h35,
8'h65,
8'h65,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'he5,
8'h25,
8'h25,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'ha5,
8'ha5,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'hc5,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'h35,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'hd5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h65,
8'h25,
8'h15,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'ha5,
8'h95,
8'h95,
8'h55,
8'h55,
8'h55,
8'h55,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'hc5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h35,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h45,
8'h45,
8'h25,
8'h15,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'ha5,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'hc5,
8'h25,
8'h25,
8'h25,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'hf5,
8'h65,
8'h25,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'ha5,
8'h55,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'h85,
8'h85,
8'h85,
8'h85,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'h25,
8'h25,
8'hc5,
8'h35,
8'hd5,
8'h35,
8'h35,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h35,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h95,
8'h85,
8'h85,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h85,
8'h85,
8'h85,
8'h55,
8'h55,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'h25,
8'h25,
8'hc5,
8'h35,
8'h35,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h95,
8'h95,
8'h95,
8'h55,
8'h55,
8'h55,
8'h95,
8'ha5,
8'ha5,
8'h25,
8'he5,
8'h25,
8'h25,
8'h35,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h25,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'ha5,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h95,
8'h25,
8'he5,
8'he5,
8'he5,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'he5,
8'he5,
8'ha5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h45,
8'h25,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'ha5,
8'h55,
8'h55,
8'h55,
8'h55,
8'h95,
8'he5,
8'h15,
8'h15,
8'h15,
8'h15,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'he5,
8'he5,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'h15,
8'he5,
8'he5,
8'ha5,
8'ha5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h45,
8'h45,
8'h25,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h95,
8'h55,
8'h55,
8'h55,
8'h95,
8'h15,
8'h15,
8'he5,
8'h25,
8'h95,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h95,
8'h95,
8'h25,
8'h25,
8'he5,
8'h15,
8'he5,
8'h25,
8'ha5,
8'h95,
8'ha5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h65,
8'h25,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h95,
8'h55,
8'h55,
8'h55,
8'h15,
8'h15,
8'h25,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h95,
8'h55,
8'h55,
8'h95,
8'h95,
8'h95,
8'ha5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h55,
8'h55,
8'h55,
8'h25,
8'h15,
8'h25,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h95,
8'h55,
8'h55,
8'he5,
8'h15,
8'h95,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h55,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h25,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h95,
8'h55,
8'h55,
8'h15,
8'h15,
8'h95,
8'h55,
8'h55,
8'h55,
8'h55,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'h95,
8'ha5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h45,
8'h25,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h95,
8'h55,
8'h95,
8'he5,
8'h25,
8'ha5,
8'h95,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'ha5,
8'h95,
8'ha5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h45,
8'h25,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'ha5,
8'ha5,
8'ha5,
8'h25,
8'h25,
8'ha5,
8'ha5,
8'ha5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'ha5,
8'ha5,
8'hd5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h65,
8'h65,
8'hc5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'hd5,
8'ha5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'hc5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hc5,
8'hc5,
8'h25,
8'h25,
8'h25,
8'h35,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'hc5,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'hc5,
8'h25,
8'hc5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hc5,
8'h25,
8'hc5,
8'h25,
8'hc5,
8'hd5,
8'h35,
8'h25,
8'hc5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h25,
8'h25,
8'h35,
8'h35,
8'hd5,
8'hc5,
8'hc5,
8'h35,
8'hd5,
8'h25,
8'hc5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'hc5,
8'hc5,
8'hc5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'h25,
8'hc5,
8'h35,
8'h35,
8'h35,
8'hc5,
8'h25,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'hc5,
8'h35,
8'h35,
8'h35,
8'h25,
8'hc5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'h35,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'hc5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h35,
8'h25,
8'h25,
8'hd5,
8'h35,
8'hd5,
8'h25,
8'hc5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hc5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h25,
8'h35,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'hc5,
8'h35,
8'hd5,
8'h35,
8'h25,
8'h25,
8'hc5,
8'h35,
8'h35,
8'h35,
8'hd5,
8'h35,
8'h35,
8'h25,
8'h25,
8'h25,
8'h25,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h35,
8'h35,
8'h35,
8'hd5,
8'h25,
8'hc5,
8'hd5,
8'h35,
8'h35,
8'hd5,
8'hc5,
8'hc5,
8'h35,
8'h35,
8'h35,
8'h35,
8'hc5,
8'hc5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h35,
8'hd5,
8'h35,
8'h35,
8'h25,
8'hc5,
8'h35,
8'h25,
8'h35,
8'h35,
8'hd5,
8'h25,
8'hc5,
8'h25,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'he5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'hc5,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'h35,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'hc5,
8'h25,
8'h35,
8'h35,
8'h35,
8'hc5,
8'hc5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hc5,
8'hc5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'hd5,
8'h35,
8'hd5,
8'h25,
8'h25,
8'hd5,
8'hc5,
8'h25,
8'h35,
8'h35,
8'h35,
8'h25,
8'hc5,
8'hc5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'hc5,
8'hc5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hc5,
8'h25,
8'hc5,
8'hc5,
8'h35,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'h25,
8'hc5,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'hd5,
8'h35,
8'h35,
8'h25,
8'h25,
8'h25,
8'h25,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'h25,
8'hc5,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h25,
8'h25,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'hd5,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'h35,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'h25,
8'h25,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'h25,
8'h25,
8'h25,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'h35,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hd5,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'hc5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'hc5,
8'hc5,
8'hc5,
8'hc5,
8'h35,
8'h35,
8'h35,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'hc5,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h25,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h05,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'hd4,
8'hc4,
8'h24,
8'h24,
8'hc4,
8'h24,
8'he4,
8'he4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h24,
8'h24,
8'h24,
8'hc4,
8'h34,
8'h24,
8'h24,
8'hc4,
8'h34,
8'h24,
8'h14,
8'h14,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h34,
8'hd4,
8'hd4,
8'h34,
8'hd4,
8'hc4,
8'h14,
8'h14,
8'he4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hc4,
8'h14,
8'h14,
8'he4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hc4,
8'h14,
8'h14,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h64,
8'h64,
8'h64,
8'h34,
8'hd4,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hc4,
8'he4,
8'he4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'hf4,
8'h44,
8'h64,
8'h34,
8'hc4,
8'hc4,
8'h34,
8'h24,
8'he4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'hc4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hc4,
8'he4,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'h44,
8'h44,
8'h64,
8'h34,
8'h34,
8'hc4,
8'h34,
8'h34,
8'hd4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h04,
8'h24,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h24,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h34,
8'h44,
8'h44,
8'h64,
8'h34,
8'h34,
8'hc4,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'h34,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h64,
8'h64,
8'h34,
8'hc4,
8'hc4,
8'h34,
8'h34,
8'h34,
8'hd4,
8'h34,
8'h34,
8'hc4,
8'h24,
8'h24,
8'h24,
8'hc4,
8'hc4,
8'hd4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h24,
8'h04,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'hd4,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'h34,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'hc4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'ha4,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'h24,
8'he4,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'h34,
8'h24,
8'h24,
8'h24,
8'h24,
8'hc4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'ha4,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'h14,
8'h24,
8'h44,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'h34,
8'h34,
8'h34,
8'hd4,
8'h34,
8'h24,
8'h24,
8'h24,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'ha4,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'h14,
8'h24,
8'h44,
8'h44,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'h34,
8'h34,
8'hd4,
8'h34,
8'hc4,
8'h24,
8'h24,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h84,
8'h84,
8'h84,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'h54,
8'ha4,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'h14,
8'h24,
8'h64,
8'hf4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h34,
8'h34,
8'hc4,
8'h24,
8'h24,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h54,
8'h54,
8'h54,
8'h84,
8'h84,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h84,
8'h94,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'h34,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h34,
8'h24,
8'h24,
8'he4,
8'h24,
8'ha4,
8'ha4,
8'h94,
8'h54,
8'h54,
8'h54,
8'h94,
8'h24,
8'h94,
8'h94,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'ha4,
8'he4,
8'he4,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'he4,
8'he4,
8'h24,
8'h94,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'ha4,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'ha4,
8'ha4,
8'he4,
8'he4,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'h14,
8'he4,
8'he4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'h14,
8'h14,
8'h14,
8'h14,
8'he4,
8'h94,
8'h54,
8'h54,
8'h54,
8'h54,
8'ha4,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h44,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'ha4,
8'h94,
8'ha4,
8'h24,
8'he4,
8'he4,
8'he4,
8'h24,
8'h24,
8'h94,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h94,
8'h24,
8'he4,
8'h14,
8'h14,
8'h94,
8'h54,
8'h54,
8'h54,
8'h94,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h44,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h94,
8'h14,
8'h14,
8'h54,
8'h54,
8'h54,
8'h94,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h64,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h24,
8'h14,
8'h24,
8'h54,
8'h54,
8'h94,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h54,
8'h94,
8'h14,
8'he4,
8'h54,
8'h54,
8'h94,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'h94,
8'h94,
8'h94,
8'h94,
8'h54,
8'h54,
8'h54,
8'h94,
8'h14,
8'h14,
8'h54,
8'h54,
8'h94,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'h24,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'ha4,
8'h94,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'ha4,
8'h94,
8'ha4,
8'h24,
8'he4,
8'h94,
8'h54,
8'ha4,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'h24,
8'h44,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hd4,
8'ha4,
8'ha4,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h94,
8'ha4,
8'ha4,
8'h24,
8'h24,
8'ha4,
8'ha4,
8'ha4,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'h64,
8'h44,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h34,
8'h24,
8'h24,
8'hc4,
8'hc4,
8'hc4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'hc4,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'ha4,
8'hd4,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'h64,
8'h64,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'hc4,
8'h24,
8'hc4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h64,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'hc4,
8'h24,
8'h34,
8'hd4,
8'hc4,
8'hc4,
8'hc4,
8'h24,
8'hc4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'hc4,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hc4,
8'h24,
8'hd4,
8'h34,
8'hc4,
8'hc4,
8'hd4,
8'h34,
8'h34,
8'hc4,
8'h24,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hc4,
8'h24,
8'h34,
8'h34,
8'h34,
8'hc4,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'h24,
8'hc4,
8'h34,
8'h34,
8'h34,
8'hc4,
8'h24,
8'hc4,
8'h24,
8'he4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'hc4,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h34,
8'h24,
8'h34,
8'h34,
8'h34,
8'h34,
8'hc4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hc4,
8'h24,
8'h34,
8'h34,
8'hd4,
8'h24,
8'h24,
8'h34,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'hc4,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hc4,
8'hc4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h24,
8'hd4,
8'h34,
8'h34,
8'hd4,
8'hc4,
8'h24,
8'h34,
8'h34,
8'h34,
8'h34,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h24,
8'h24,
8'h24,
8'hc4,
8'h34,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h24,
8'h24,
8'h24,
8'h34,
8'hd4,
8'h34,
8'h34,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'hc4,
8'hc4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'hc4,
8'h24,
8'hc4,
8'h34,
8'h34,
8'h24,
8'hc4,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'h34,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'hc4,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'he4,
8'h24,
8'h24,
8'h24,
8'hd4,
8'h34,
8'h34,
8'h24,
8'h34,
8'hc4,
8'h24,
8'h34,
8'h34,
8'hd4,
8'h34,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h34,
8'h24,
8'h34,
8'h34,
8'hd4,
8'h34,
8'h34,
8'hd4,
8'h34,
8'hc4,
8'hc4,
8'h24,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hc4,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'hc4,
8'hc4,
8'hc4,
8'h34,
8'h34,
8'h34,
8'h24,
8'hc4,
8'hd4,
8'h24,
8'h24,
8'hd4,
8'h34,
8'h34,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'hc4,
8'h24,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h24,
8'h24,
8'h24,
8'hc4,
8'h34,
8'h34,
8'hd4,
8'h24,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h34,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'h24,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'hc4,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'hd4,
8'hd4,
8'hd4,
8'hd4,
8'h34,
8'h24,
8'hc4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h34,
8'h34,
8'h34,
8'hc4,
8'hc4,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'hc4,
8'h24,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'h24,
8'hd4,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04,
8'h04

	};


	
	    
 always_comb begin:tank_select
 
 case(tankSelection)
 
 2'b00: begin
  data = R_ROM[addr + 3500 * Direction];
 
 end
 
 2'b01: begin
  data = Y_ROM[addr + 3500 * Direction]; 
 end
 
 2'b10: begin
  data = B_ROM[addr + 3500 * Direction];
 end
 
 2'b11: begin
  data = B_ROM[addr + 3500 * Direction];
 end
 
 default:;
 
 endcase
 
 end



endmodule  






