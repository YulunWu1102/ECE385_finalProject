module gameover_rom ( input [12:0]	addr,
						output [3:0]	data
					 );

				
	// ROM definition
// 150 x 50				
	parameter [0:7499][3:0] ROM = {

4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h3,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h3,
4'h3,
4'h3,
4'hd,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h3,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h3,
4'h3,
4'hd,
4'hd,
4'hc,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'hd,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h3,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h2,
4'he,
4'h1,
4'he,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'hd,
4'hd,
4'hd,
4'h2,
4'h2,
4'h1,
4'h1,
4'h2,
4'he,
4'h1,
4'he,
4'h2,
4'h2,
4'hd,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'hc,
4'hd,
4'h2,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h2,
4'h1,
4'h1,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'he,
4'h1,
4'he,
4'h2,
4'h2,
4'hd,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h3,
4'h2,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'he,
4'h1,
4'he,
4'h2,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h3,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'hc,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h3,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'h2,
4'hd,
4'h3,
4'hc,
4'he,
4'h1,
4'h1,
4'h1,
4'h3,
4'h2,
4'h1,
4'h1,
4'h1,
4'he,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hc,
4'h2,
4'he,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'h3,
4'h2,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'he,
4'he,
4'he,
4'he,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hc,
4'h1,
4'h1,
4'h1,
4'he,
4'hc,
4'he,
4'h1,
4'h2,
4'hc,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hc,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'he,
4'he,
4'he,
4'he,
4'h1,
4'he,
4'h3,
4'hc,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'he,
4'he,
4'h1,
4'h2,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hc,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'h2,
4'he,
4'hc,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'h3,
4'he,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hc,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'he,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'hc,
4'hd,
4'hd,
4'hd,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hc,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'hc,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h2,
4'he,
4'h1,
4'he,
4'he,
4'he,
4'he,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h2,
4'hc,
4'h1,
4'h1,
4'h1,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'he,
4'h1,
4'h1,
4'h1,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h2,
4'he,
4'h1,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'h1,
4'he,
4'hc,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'h3,
4'h2,
4'h2,
4'h1,
4'he,
4'h2,
4'h3,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'h1,
4'h1,
4'h1,
4'h1,
4'hd,
4'hd,
4'h2,
4'h2,
4'h1,
4'h1,
4'h1,
4'h1,
4'he,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'h2,
4'hd,
4'h2,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'he,
4'he,
4'he,
4'hc,
4'h3,
4'he,
4'he,
4'he,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'he,
4'he,
4'he,
4'hd,
4'h2,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hc,
4'he,
4'h2,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'h2,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'he,
4'he,
4'he,
4'he,
4'hd,
4'hd,
4'hd,
4'hc,
4'he,
4'he,
4'he,
4'he,
4'he,
4'hc,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd,
4'hd


        };

	assign data = ROM[addr];

endmodule 