module rtank_rom ( input [15:0]	addr,
						output [3:0]	data
					 );

	parameter ADDR_WIDTH = 16;
   parameter DATA_WIDTH =  4;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {


<<<<<<< HEAD
4'h9,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h2,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h1,
4'h1,
4'h1,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h3,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
=======



4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h2
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h1
4'h1
4'h1
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h3
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
4'h0
>>>>>>> f4970183a89d1e33ee5e7378306e7847bbad6afa

// above are rtank



        };

	assign data = ROM[addr];

endmodule  