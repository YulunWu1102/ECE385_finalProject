module exp_rom ( input [13:0]	addr,						 
						 output [4:0]	data
					 );

	parameter ADDR_WIDTH = 9;
   parameter DATA_WIDTH =  4;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition
	//20 x 20 explosion

		

	parameter [0:399][3:0] EXP = {
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h7,
4'h0,
4'h0,
4'h0,
4'h0,
4'h7,
4'h0,
4'h0,
4'h0,
4'h0,
4'h7,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h7,
4'h7,
4'h7,
4'h0,
4'h0,
4'hb,
4'h4,
4'h0,
4'h7,
4'h7,
4'h7,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h7,
4'h7,
4'h7,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h7,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h4,
4'h4,
4'h4,
4'hb,
4'h4,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h4,
4'hb,
4'hb,
4'hb,
4'hb,
4'h7,
4'h4,
4'h6,
4'h4,
4'h4,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'hf,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'hb,
4'hb,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h4,
4'h4,
4'hb,
4'hb,
4'h4,
4'h4,
4'h4,
4'hb,
4'hb,
4'hf,
4'h4,
4'h4,
4'hb,
4'h7,
4'he,
4'h0,
4'h0,
4'h0,
4'h7,
4'h7,
4'h4,
4'h4,
4'hb,
4'hb,
4'h4,
4'h6,
4'h4,
4'h4,
4'hb,
4'h4,
4'h4,
4'h4,
4'hb,
4'h7,
4'h0,
4'h0,
4'h0,
4'h7,
4'h7,
4'h7,
4'hb,
4'h4,
4'h4,
4'hb,
4'h7,
4'hb,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h2,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h6,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'h4,
4'hb,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h4,
4'hb,
4'h4,
4'h4,
4'h4,
4'h4,
4'h7,
4'h7,
4'h7,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h7,
4'h7,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h7,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h7,
4'h4,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'he,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0,
4'h0

	};

	assign data = EXP[addr];

endmodule  